module clock(AM,A,B);
input A,B;
output AM;
assign AM = A;
endmodule